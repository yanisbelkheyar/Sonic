--------------------------------------------------------------------------------
--! @file       sonic512_pkg.vhd
--! @brief      Package for the sonic512 permutation.
--!
--! @author     
--------------------------------------------------------------------------------

library IEEE;
    use IEEE.std_logic_1164.all;

library work;

package sonic512_pkg is
    
	-- reset
	constant active_rst : std_logic := '0';
	
    -- size
    constant SIZE         : integer := 512;
    -- number of rounds
    constant nrRounds     : integer := 16;
    
    --types
    type rc_state is array(integer range 0 to (nrRounds - 1)) of std_logic_vector(0 to SIZE/2-1);
    type state is array(integer range 0 to (nrRounds - 1)) of std_logic_vector(0 to SIZE-1);
    type offsets is array(integer range 0 to (nrRounds - 1)) of integer;
    
    constant round_constants : rc_state := (x"8000000080000000800000008000000080000000800000000000000000000000",  -- f9
                                            x"8000000080000000800000000000000000000000000000008000000000000000",  -- 47
                                            x"8000000080000000800000008000000000000000800000000000000080000000",  -- eb
                                            x"8000000080000000800000000000000080000000800000000000000000000000",  -- 37
                                            x"8000000000000000800000008000000000000000800000000000000000000000",  -- 69
                                            x"8000000080000000000000008000000080000000800000000000000000000000",  -- 3b
                                            x"8000000000000000800000000000000000000000800000000000000000000000",  -- 49
                                            x"0000000080000000000000008000000080000000800000000000000000000000",  -- 3a
                                            x"0000000080000000000000008000000080000000000000000000000000000000",  -- b0
                                            x"8000000000000000800000008000000080000000800000008000000000000000",  -- 7d
                                            x"8000000000000000800000000000000080000000800000000000000080000000",  -- 5b
                                            x"0000000080000000000000008000000000000000000000008000000000000000",  -- 4a
                                            x"0000000000000000000000008000000080000000000000000000000080000000",  -- 32
                                            x"8000000000000000000000000000000080000000800000008000000000000000",  -- 71
                                            x"8000000000000000800000008000000080000000800000000000000080000000",  -- 7b
                                            x"8000000080000000000000008000000000000000000000008000000000000000"); -- 4b
    
    constant pi_1_offsets : offsets := (239,33,207,65,175,97,143,129,111,161,79,193,47,225,15,1);
    constant pi_5_offsets : offsets := (171,165,11,69,107,229,203,133,43,37,139,197,235,101,75,5);
    constant pi_7_offsets : offsets := (137,231,169,199,201,167,233,135,9,103,41,71,73,39,105,7);
    constant pi_32_offsets : offsets := (224,32,224,32,224,32,224,32,224,32,224,32,224,32,224,32);
	
    
end package;

